library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

library work;
use work.FRAME_PACK.all;

entity CRC32_GEN is
	port(
		CLK, RST : in std_logic;
		
		INPUT : in std_logic_vector(7 downto 0);
		N : in integer;
		OUTPUT : out std_logic_vector(31 downto 0)
	);
end CRC32_GEN;

architecture behavioral of CRC32_GEN is
signal CRC32_LUT : CRC32_ARR;
begin
p_decode:process(CLK) is
constant CRC32_POLY : std_logic_vector(31 downto 0) := x"04C11DB7";
variable CRC32 : std_logic_vector(31 downto 0);
variable i : integer;
variable ref_byte : std_logic_vector(7 downto 0);
variable LUT_search : std_logic_vector(7 downto 0);
begin
if(rising_edge(CLK)) then
	if(RST = '1') then
		i := 0;	
		CRC32 := (others => '1'); -- initial CRC
	else
		if(i < N) then
			-- reflect the input data
			for k in 0 to 7 loop
				ref_byte(k) := INPUT(7 - k);
			end loop;
			LUT_search := (CRC32(31 downto 24) AND x"FF") XOR ref_byte;
			CRC32 := (CRC32(23 downto 0) & x"00") XOR CRC32_LUT(to_integer(unsigned(LUT_search)));
			i := i + 1;
		else
			for k in 0 to 31 loop
				OUTPUT(k) <= CRC32(31-k) XOR '1';
			end loop;
		end if;
	end if;
end if;
end process;

CRC32_LUT(0) <= x"00000000";
CRC32_LUT(1) <= x"04C11DB7";
CRC32_LUT(2) <= x"09823B6E";
CRC32_LUT(3) <= x"0D4326D9";
CRC32_LUT(4) <= x"130476DC";
CRC32_LUT(5) <= x"17C56B6B";
CRC32_LUT(6) <= x"1A864DB2";
CRC32_LUT(7) <= x"1E475005";
CRC32_LUT(8) <= x"2608EDB8";
CRC32_LUT(9) <= x"22C9F00F";
CRC32_LUT(10) <= x"2F8AD6D6";
CRC32_LUT(11) <= x"2B4BCB61";
CRC32_LUT(12) <= x"350C9B64";
CRC32_LUT(13) <= x"31CD86D3";
CRC32_LUT(14) <= x"3C8EA00A";
CRC32_LUT(15) <= x"384FBDBD";
CRC32_LUT(16) <= x"4C11DB70";
CRC32_LUT(17) <= x"48D0C6C7";
CRC32_LUT(18) <= x"4593E01E";
CRC32_LUT(19) <= x"4152FDA9";
CRC32_LUT(20) <= x"5F15ADAC";
CRC32_LUT(21) <= x"5BD4B01B";
CRC32_LUT(22) <= x"569796C2";
CRC32_LUT(23) <= x"52568B75";
CRC32_LUT(24) <= x"6A1936C8";
CRC32_LUT(25) <= x"6ED82B7F";
CRC32_LUT(26) <= x"639B0DA6";
CRC32_LUT(27) <= x"675A1011";
CRC32_LUT(28) <= x"791D4014";
CRC32_LUT(29) <= x"7DDC5DA3";
CRC32_LUT(30) <= x"709F7B7A";
CRC32_LUT(31) <= x"745E66CD";
CRC32_LUT(32) <= x"9823B6E0";
CRC32_LUT(33) <= x"9CE2AB57";
CRC32_LUT(34) <= x"91A18D8E";
CRC32_LUT(35) <= x"95609039";
CRC32_LUT(36) <= x"8B27C03C";
CRC32_LUT(37) <= x"8FE6DD8B";
CRC32_LUT(38) <= x"82A5FB52";
CRC32_LUT(39) <= x"8664E6E5";
CRC32_LUT(40) <= x"BE2B5B58";
CRC32_LUT(41) <= x"BAEA46EF";
CRC32_LUT(42) <= x"B7A96036";
CRC32_LUT(43) <= x"B3687D81";
CRC32_LUT(44) <= x"AD2F2D84";
CRC32_LUT(45) <= x"A9EE3033";
CRC32_LUT(46) <= x"A4AD16EA";
CRC32_LUT(47) <= x"A06C0B5D";
CRC32_LUT(48) <= x"D4326D90";
CRC32_LUT(49) <= x"D0F37027";
CRC32_LUT(50) <= x"DDB056FE";
CRC32_LUT(51) <= x"D9714B49";
CRC32_LUT(52) <= x"C7361B4C";
CRC32_LUT(53) <= x"C3F706FB";
CRC32_LUT(54) <= x"CEB42022";
CRC32_LUT(55) <= x"CA753D95";
CRC32_LUT(56) <= x"F23A8028";
CRC32_LUT(57) <= x"F6FB9D9F";
CRC32_LUT(58) <= x"FBB8BB46";
CRC32_LUT(59) <= x"FF79A6F1";
CRC32_LUT(60) <= x"E13EF6F4";
CRC32_LUT(61) <= x"E5FFEB43";
CRC32_LUT(62) <= x"E8BCCD9A";
CRC32_LUT(63) <= x"EC7DD02D";
CRC32_LUT(64) <= x"34867077";
CRC32_LUT(65) <= x"30476DC0";
CRC32_LUT(66) <= x"3D044B19";
CRC32_LUT(67) <= x"39C556AE";
CRC32_LUT(68) <= x"278206AB";
CRC32_LUT(69) <= x"23431B1C";
CRC32_LUT(70) <= x"2E003DC5";
CRC32_LUT(71) <= x"2AC12072";
CRC32_LUT(72) <= x"128E9DCF";
CRC32_LUT(73) <= x"164F8078";
CRC32_LUT(74) <= x"1B0CA6A1";
CRC32_LUT(75) <= x"1FCDBB16";
CRC32_LUT(76) <= x"018AEB13";
CRC32_LUT(77) <= x"054BF6A4";
CRC32_LUT(78) <= x"0808D07D";
CRC32_LUT(79) <= x"0CC9CDCA";
CRC32_LUT(80) <= x"7897AB07";
CRC32_LUT(81) <= x"7C56B6B0";
CRC32_LUT(82) <= x"71159069";
CRC32_LUT(83) <= x"75D48DDE";
CRC32_LUT(84) <= x"6B93DDDB";
CRC32_LUT(85) <= x"6F52C06C";
CRC32_LUT(86) <= x"6211E6B5";
CRC32_LUT(87) <= x"66D0FB02";
CRC32_LUT(88) <= x"5E9F46BF";
CRC32_LUT(89) <= x"5A5E5B08";
CRC32_LUT(90) <= x"571D7DD1";
CRC32_LUT(91) <= x"53DC6066";
CRC32_LUT(92) <= x"4D9B3063";
CRC32_LUT(93) <= x"495A2DD4";
CRC32_LUT(94) <= x"44190B0D";
CRC32_LUT(95) <= x"40D816BA";
CRC32_LUT(96) <= x"ACA5C697";
CRC32_LUT(97) <= x"A864DB20";
CRC32_LUT(98) <= x"A527FDF9";
CRC32_LUT(99) <= x"A1E6E04E";
CRC32_LUT(100) <= x"BFA1B04B";
CRC32_LUT(101) <= x"BB60ADFC";
CRC32_LUT(102) <= x"B6238B25";
CRC32_LUT(103) <= x"B2E29692";
CRC32_LUT(104) <= x"8AAD2B2F";
CRC32_LUT(105) <= x"8E6C3698";
CRC32_LUT(106) <= x"832F1041";
CRC32_LUT(107) <= x"87EE0DF6";
CRC32_LUT(108) <= x"99A95DF3";
CRC32_LUT(109) <= x"9D684044";
CRC32_LUT(110) <= x"902B669D";
CRC32_LUT(111) <= x"94EA7B2A";
CRC32_LUT(112) <= x"E0B41DE7";
CRC32_LUT(113) <= x"E4750050";
CRC32_LUT(114) <= x"E9362689";
CRC32_LUT(115) <= x"EDF73B3E";
CRC32_LUT(116) <= x"F3B06B3B";
CRC32_LUT(117) <= x"F771768C";
CRC32_LUT(118) <= x"FA325055";
CRC32_LUT(119) <= x"FEF34DE2";
CRC32_LUT(120) <= x"C6BCF05F";
CRC32_LUT(121) <= x"C27DEDE8";
CRC32_LUT(122) <= x"CF3ECB31";
CRC32_LUT(123) <= x"CBFFD686";
CRC32_LUT(124) <= x"D5B88683";
CRC32_LUT(125) <= x"D1799B34";
CRC32_LUT(126) <= x"DC3ABDED";
CRC32_LUT(127) <= x"D8FBA05A";
CRC32_LUT(128) <= x"690CE0EE";
CRC32_LUT(129) <= x"6DCDFD59";
CRC32_LUT(130) <= x"608EDB80";
CRC32_LUT(131) <= x"644FC637";
CRC32_LUT(132) <= x"7A089632";
CRC32_LUT(133) <= x"7EC98B85";
CRC32_LUT(134) <= x"738AAD5C";
CRC32_LUT(135) <= x"774BB0EB";
CRC32_LUT(136) <= x"4F040D56";
CRC32_LUT(137) <= x"4BC510E1";
CRC32_LUT(138) <= x"46863638";
CRC32_LUT(139) <= x"42472B8F";
CRC32_LUT(140) <= x"5C007B8A";
CRC32_LUT(141) <= x"58C1663D";
CRC32_LUT(142) <= x"558240E4";
CRC32_LUT(143) <= x"51435D53";
CRC32_LUT(144) <= x"251D3B9E";
CRC32_LUT(145) <= x"21DC2629";
CRC32_LUT(146) <= x"2C9F00F0";
CRC32_LUT(147) <= x"285E1D47";
CRC32_LUT(148) <= x"36194D42";
CRC32_LUT(149) <= x"32D850F5";
CRC32_LUT(150) <= x"3F9B762C";
CRC32_LUT(151) <= x"3B5A6B9B";
CRC32_LUT(152) <= x"0315D626";
CRC32_LUT(153) <= x"07D4CB91";
CRC32_LUT(154) <= x"0A97ED48";
CRC32_LUT(155) <= x"0E56F0FF";
CRC32_LUT(156) <= x"1011A0FA";
CRC32_LUT(157) <= x"14D0BD4D";
CRC32_LUT(158) <= x"19939B94";
CRC32_LUT(159) <= x"1D528623";
CRC32_LUT(160) <= x"F12F560E";
CRC32_LUT(161) <= x"F5EE4BB9";
CRC32_LUT(162) <= x"F8AD6D60";
CRC32_LUT(163) <= x"FC6C70D7";
CRC32_LUT(164) <= x"E22B20D2";
CRC32_LUT(165) <= x"E6EA3D65";
CRC32_LUT(166) <= x"EBA91BBC";
CRC32_LUT(167) <= x"EF68060B";
CRC32_LUT(168) <= x"D727BBB6";
CRC32_LUT(169) <= x"D3E6A601";
CRC32_LUT(170) <= x"DEA580D8";
CRC32_LUT(171) <= x"DA649D6F";
CRC32_LUT(172) <= x"C423CD6A";
CRC32_LUT(173) <= x"C0E2D0DD";
CRC32_LUT(174) <= x"CDA1F604";
CRC32_LUT(175) <= x"C960EBB3";
CRC32_LUT(176) <= x"BD3E8D7E";
CRC32_LUT(177) <= x"B9FF90C9";
CRC32_LUT(178) <= x"B4BCB610";
CRC32_LUT(179) <= x"B07DABA7";
CRC32_LUT(180) <= x"AE3AFBA2";
CRC32_LUT(181) <= x"AAFBE615";
CRC32_LUT(182) <= x"A7B8C0CC";
CRC32_LUT(183) <= x"A379DD7B";
CRC32_LUT(184) <= x"9B3660C6";
CRC32_LUT(185) <= x"9FF77D71";
CRC32_LUT(186) <= x"92B45BA8";
CRC32_LUT(187) <= x"9675461F";
CRC32_LUT(188) <= x"8832161A";
CRC32_LUT(189) <= x"8CF30BAD";
CRC32_LUT(190) <= x"81B02D74";
CRC32_LUT(191) <= x"857130C3";
CRC32_LUT(192) <= x"5D8A9099";
CRC32_LUT(193) <= x"594B8D2E";
CRC32_LUT(194) <= x"5408ABF7";
CRC32_LUT(195) <= x"50C9B640";
CRC32_LUT(196) <= x"4E8EE645";
CRC32_LUT(197) <= x"4A4FFBF2";
CRC32_LUT(198) <= x"470CDD2B";
CRC32_LUT(199) <= x"43CDC09C";
CRC32_LUT(200) <= x"7B827D21";
CRC32_LUT(201) <= x"7F436096";
CRC32_LUT(202) <= x"7200464F";
CRC32_LUT(203) <= x"76C15BF8";
CRC32_LUT(204) <= x"68860BFD";
CRC32_LUT(205) <= x"6C47164A";
CRC32_LUT(206) <= x"61043093";
CRC32_LUT(207) <= x"65C52D24";
CRC32_LUT(208) <= x"119B4BE9";
CRC32_LUT(209) <= x"155A565E";
CRC32_LUT(210) <= x"18197087";
CRC32_LUT(211) <= x"1CD86D30";
CRC32_LUT(212) <= x"029F3D35";
CRC32_LUT(213) <= x"065E2082";
CRC32_LUT(214) <= x"0B1D065B";
CRC32_LUT(215) <= x"0FDC1BEC";
CRC32_LUT(216) <= x"3793A651";
CRC32_LUT(217) <= x"3352BBE6";
CRC32_LUT(218) <= x"3E119D3F";
CRC32_LUT(219) <= x"3AD08088";
CRC32_LUT(220) <= x"2497D08D";
CRC32_LUT(221) <= x"2056CD3A";
CRC32_LUT(222) <= x"2D15EBE3";
CRC32_LUT(223) <= x"29D4F654";
CRC32_LUT(224) <= x"C5A92679";
CRC32_LUT(225) <= x"C1683BCE";
CRC32_LUT(226) <= x"CC2B1D17";
CRC32_LUT(227) <= x"C8EA00A0";
CRC32_LUT(228) <= x"D6AD50A5";
CRC32_LUT(229) <= x"D26C4D12";
CRC32_LUT(230) <= x"DF2F6BCB";
CRC32_LUT(231) <= x"DBEE767C";
CRC32_LUT(232) <= x"E3A1CBC1";
CRC32_LUT(233) <= x"E760D676";
CRC32_LUT(234) <= x"EA23F0AF";
CRC32_LUT(235) <= x"EEE2ED18";
CRC32_LUT(236) <= x"F0A5BD1D";
CRC32_LUT(237) <= x"F464A0AA";
CRC32_LUT(238) <= x"F9278673";
CRC32_LUT(239) <= x"FDE69BC4";
CRC32_LUT(240) <= x"89B8FD09";
CRC32_LUT(241) <= x"8D79E0BE";
CRC32_LUT(242) <= x"803AC667";
CRC32_LUT(243) <= x"84FBDBD0";
CRC32_LUT(244) <= x"9ABC8BD5";
CRC32_LUT(245) <= x"9E7D9662";
CRC32_LUT(246) <= x"933EB0BB";
CRC32_LUT(247) <= x"97FFAD0C";
CRC32_LUT(248) <= x"AFB010B1";
CRC32_LUT(249) <= x"AB710D06";
CRC32_LUT(250) <= x"A6322BDF";
CRC32_LUT(251) <= x"A2F33668";
CRC32_LUT(252) <= x"BCB4666D";
CRC32_LUT(253) <= x"B8757BDA";
CRC32_LUT(254) <= x"B5365D03";
CRC32_LUT(255) <= x"B1F740B4";
end behavioral;
